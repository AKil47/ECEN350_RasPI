`timescale 1ns / 1ps

`define OPCODE_MOVZ   9'b110100101
`define OPCODE_ORRREG 11'b00101010000
`define OPCODE_STUR   11'b11111000000
`define OPCODE_LDUR   11'b11111000010

/*
 * Module: InstructionMemory
 *
 * Implements read-only instruction memory
 * 
 */
module InstructionMemory(Data, Address);
   parameter T_rd = 20;
   parameter MemSize = 40;
   
   output [31:0] Data;
   input [63:0]  Address;
   reg [31:0] 	 Data;
   
   /*
    * ECEN 350 Processor Test Functions
    * Texas A&M University
    */
    
    reg [31:0] test;
    
    

   
   always @ (Address) begin

      case(Address)

	/* Test Program 1:
	 * Program loads constants from the data memory. Uses these constants to test
	 * the following instructions: LDUR, ORR, AND, CBZ, ADD, SUB, STUR and B.
	 * 
	 * Assembly code for test:
	 * 
	 * 0: LDUR X9, [XZR, 0x0]    //Load 1 into x9
	 * 4: LDUR X10, [XZR, 0x8]   //Load a into x10
	 * 8: LDUR X11, [XZR, 0x10]  //Load 5 into x11
	 * C: LDUR X12, [XZR, 0x18]  //Load big constant into x12
	 * 10: LDUR X13, [XZR, 0x20]  //load a 0 into X13
	 * 
	 * 14: ORR X10, X10, X11  //Create mask of 0xf
	 * 18: AND X12, X12, X10  //Mask off low order bits of big constant
	 * 
	 * loop:
	 * 1C: CBZ X12, end  //while X12 is not 0
	 * 20: ADD X13, X13, X9  //Increment counter in X13
	 * 24: SUB X12, X12, X9  //Decrement remainder of big constant in X12
	 * 28: B loop  //Repeat till X12 is 0
	 * 2C: STUR X13, [XZR, 0x20]  //store back the counter value into the memory location 0x20
	 */
	

	63'h000: Data = 32'hf84003e9;
	63'h004: Data = 32'hf84083ea;
	63'h008: Data = 32'hf84103eb;
	63'h00c: Data = 32'hf84183ec;
	63'h010: Data = 32'hf84203ed;
	63'h014: Data = 32'haa0b014a;
	63'h018: Data = 32'h8a0a018c;
	63'h01c: Data = 32'hb400008c;
	63'h020: Data = 32'h8b0901ad;
	63'h024: Data = 32'hcb09018c;
	63'h028: Data = 32'h17fffffd;
	63'h02c: Data = 32'hf80203ed;
	63'h030: Data = 32'hf84203ed;  //One last load to place stored value on memdbus for test checking
	
	63'h034: Data = {`OPCODE_MOVZ, 2'b11, 16'h1234, 5'd9}; //MOVZ 0xh1234 LSL 48 11010010 (11 11) 0xh1234 9
	63'h038: Data = {`OPCODE_MOVZ, 2'b10, 16'h5678, 5'd10}; //MOVK 0xh5678 LSL 32              10
	63'h03c: Data = {`OPCODE_MOVZ, 2'b01, 16'h9abc, 5'd11}; //MOVK 0xh9abc LSL 16            01
	63'h040: Data = {`OPCODE_MOVZ, 2'b00, 16'hdef0, 5'd12}; //MOVK 0xhdef0
	
	63'h044: Data = {`OPCODE_ORRREG, 5'd9, 6'd0, 5'd10, 5'd9}; // OR X9 X9 X10
	63'h048: Data = {`OPCODE_ORRREG, 5'd9, 6'd0, 5'd11, 5'd9}; // OR X9 X9 X10
	63'h04c: Data = {`OPCODE_ORRREG, 5'd9, 6'd0, 5'd12, 5'd9}; // OR X9 X9 X10
	
	63'h050: Data = {`OPCODE_STUR, 9'h28, 2'd0, 5'd31, 5'd9}; // STUR X9, [XZR, #0x28]
	63'h054: Data = {`OPCODE_LDUR, 9'h28, 2'd0, 5'd31, 5'd10}; // LDUR X10, [XZR, #0x28]	
	
	63'h058: Data = 32'hf84203ea;  //One last load to place stored value on memdbus for test checking				
					

	/* Add code for your tests here */

	
	default: Data = 32'hXXXXXXXX;
      endcase
   end
endmodule
